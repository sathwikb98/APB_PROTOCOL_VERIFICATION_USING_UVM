`define ADDR_WIDTH 9
`define DATA_WIDTH 8
`define no_of_transaction 20
